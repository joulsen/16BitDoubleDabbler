`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    22:10:55 04/28/2020 
// Design Name: 
// Module Name:    ClockedDoubleDabbler16Bit 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ClockedDoubleDabbler16Bit(
    input CLK,
    input [15:0] BIN,
    output [19:0] BCD,
    output FINISH
    );


endmodule
